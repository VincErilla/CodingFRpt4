/*
 
 Conway's Game of Life modeled in SVerilog
 
 */

module datapath ( grid, grid_evolve );

   output logic [255:0] 	grid_evolve;
   input logic [255:0] 	grid;
   
   evolve3 e0_0 (grid_evolve[0], grid[1], grid[8], grid[9], grid[0]);
   evolve5 e0_1 (grid_evolve[1], grid[0], grid[2], grid[8], grid[9], grid[10], grid[1]);
   evolve5 e0_2 (grid_evolve[2], grid[1], grid[3], grid[9], grid[10], grid[11], grid[2]);
   evolve5 e0_3 (grid_evolve[3], grid[2], grid[4], grid[10], grid[11], grid[12], grid[3]);
   evolve5 e0_4 (grid_evolve[4], grid[3], grid[5], grid[11], grid[12], grid[13], grid[4]);
   evolve5 e0_5 (grid_evolve[5], grid[4], grid[6], grid[12], grid[13], grid[14], grid[5]);
   evolve5 e0_6 (grid_evolve[6], grid[5], grid[7], grid[13], grid[14], grid[15], grid[6]);
   evolve5 e0_7 (grid_evolve[7], grid[6], grid[8], grid[14], grid[15], grid,[16], grid[7]);
   evolve5 e0_8 (grid_evolve[8], grid[7], grid[9], grid[15], grid[16], grid[17], grid[8]);
   evolve5 e0_9 (grid_evolve[9], grid[8], grid[10], grid[16], grid[17], grid[18], grid[9]);
   evolve5 e0_10 (grid_evolve[10], grid[9], grid[11], grid[17], grid[18], grid[19], grid[10]);
   evolve5 e0_11 (grid_evolve[11], grid[10], grid[12], grid[18], grid[19], grid[20], grid[11]);
   evolve5 e0_12 (grid_evolve[12], grid[11], grid[13], grid[19], grid[20], grid[21], grid[12]);
   evolve5 e0_13 (grid_evolve[13], grid[12], grid[14], grid[20], grid[21], grid[22], grid[13]);
   evolve5 e0_14 (grid_evolve[14], grid[13], grid[15], grid[21], grid[22], grid[23], grid[14]);
   evolve3 e0_15 (grid_evolve[15], grid[14], grid[22], grid[23], grid[15]);

   
   evolve5 e1_0 (grid_evolve[16], grid[0+8*1], grid[1+8*1], grid[9+8*1], grid[16+8*1], grid[17+8*1], grid[16]);
   evolve8 e1_1 (grid_evolve[17], grid[0+8*1], grid[1+8*1], grid[2+8*1], grid[8+8*1], grid[10+8*1], grid[16+8*1], grid[17+8*1], grid[18+8*1], grid[17]);
   evolve8 e1_2 (grid_evolve[18], grid[1+8*1], grid[2+8*1], grid[3+8*1], grid[9+8*1], grid[11+8*1], grid[17+8*1], grid[18+8*1], grid[19+8*1], grid[18]);
   evolve8 e1_3 (grid_evolve[19], grid[2+8*1], grid[3+8*1], grid[4+8*1], grid[10+8*1], grid[12+8*1], grid[18+8*1], grid[19+8*1], grid[20+8*1], grid[19]);
   evolve8 e1_4 (grid_evolve[20], grid[3+8*1], grid[4+8*1], grid[5+8*1], grid[11+8*1], grid[13+8*1], grid[19+8*1], grid[20+8*1], grid[21+8*1], grid[20]);
   evolve8 e1_5 (grid_evolve[21], grid[4+8*1], grid[5+8*1], grid[6+8*1], grid[12+8*1], grid[14+8*1], grid[20+8*1], grid[21+8*1], grid[22+8*1], grid[21]);
   evolve8 e1_6 (grid_evolve[22], grid[5+8*1], grid[6+8*1], grid[7+8*1], grid[13+8*1], grid[15+8*1], grid[21+8*1], grid[22+8*1], grid[23+8*1], grid[22]);
   evolve8 e1_7 (grid_evolve[23], grid[6+8*1], grid[7+8*1], grid[9+8*1], grid[14+8*1], grid[22+8*1], grid[23+8*1], grid[24+8*1], grid[23]);
   evolve8 e1_8 (grid_evolve[24], grid[15], grid[0+8*2], grid[1+8*2], grid[9+8*2], grid[31], grid[16+8*2], grid[17+8*2], grid[24]);
   evolve8 e1_9 (grid_evolve[25], grid[0+8*2], grid[1+8*2], grid[2+8*2], grid[8+8*2], grid[10+8*2], grid[16+8*2], grid[17+8*2], grid[18+8*2], grid[25]);
   evolve8 e1_10 (grid_evolve[26], grid[1+8*2], grid[2+8*2], grid[3+8*2], grid[9+8*2], grid[11+8*2], grid[17+8*2], grid[18+8*2], grid[19+8*2], grid[26]);
   evolve8 e1_11 (grid_evolve[27], grid[2+8*2], grid[3+8*2], grid[4+8*2], grid[10+8*2], grid[12+8*2], grid[18+8*2], grid[19+8*2], grid[20+8*2], grid[27]);
   evolve8 e1_12 (grid_evolve[28], grid[3+8*2], grid[4+8*2], grid[5+8*2], grid[11+8*2], grid[13+8*2], grid[19+8*2], grid[20+8*2], grid[21+8*2], grid[28]);
   evolve8 e1_13 (grid_evolve[29], grid[4+8*2], grid[5+8*2], grid[6+8*2], grid[12+8*2], grid[14+8*2], grid[20+8*2], grid[21+8*2], grid[22+8*2], grid[29]);
   evolve8 e1_14 (grid_evolve[30], grid[5+8*2], grid[6+8*2], grid[7+8*2], grid[13+8*2], grid[15+8*2], grid[21+8*2], grid[22+8*2], grid[23+8*2], grid[30]);
   evolve5 e1_15 (grid_evolve[31], grid[6+8*2], grid[7+8*2], grid[14+8*2], grid[22+8*2], grid[23+8*2], grid[31]);
 
   
   evolve5 e2_0 (grid_evolve[32], grid[0+8*3], grid[1+8*3], grid[9+8*3], grid[16+8*3], grid[17+8*3], grid[32]);
   evolve8 e2_1 (grid_evolve[33], grid[0+8*3], grid[1+8*3], grid[2+8*3], grid[8+8*3], grid[10+8*3], grid[16+8*3], grid[17+8*3], grid[18+8*3], grid[33]);
   evolve8 e2_2 (grid_evolve[34], grid[1+8*3], grid[2+8*3], grid[3+8*3], grid[9+8*3], grid[11+8*3], grid[17+8*3], grid[18+8*3], grid[19+8*3], grid[34]);
   evolve8 e2_3 (grid_evolve[35], grid[2+8*3], grid[3+8*3], grid[4+8*3], grid[10+8*3], grid[12+8*3], grid[18+8*3], grid[19+8*3], grid[20+8*3], grid[35]);
   evolve8 e2_4 (grid_evolve[36], grid[3+8*3], grid[4+8*3], grid[5+8*3], grid[11+8*3], grid[13+8*3], grid[19+8*3], grid[20+8*3], grid[21+8*3], grid[36]);
   evolve8 e2_5 (grid_evolve[37], grid[4+8*3], grid[5+8*3], grid[6+8*3], grid[12+8*3], grid[14+8*3], grid[20+8*3], grid[21+8*3], grid[22+8*3], grid[37]);
   evolve8 e2_6 (grid_evolve[38], grid[5+8*3], grid[6+8*3], grid[7+8*3], grid[13+8*3], grid[15+8*3], grid[21+8*3], grid[22+8*3], grid[23+8*3], grid[38]);
   evolve8 e2_7 (grid_evolve[39], grid[6+8*3], grid[7+8*3], grid[32], grid[14+8*3], grid[40], grid[22+8*3], grid[23+8*3], grid[48], grid[39]);  
   evolve8 e2_8 (grid_evolve[40], grid[31], grid[0+8*4], grid[1+8*4], grid[39], grid[9+8*4], grid[47], grid[16+8*4], grid[17+8*4], grid[40]);
   evolve8 e2_9 (grid_evolve[41], grid[0+8*4], grid[1+8*4], grid[2+8*4], grid[8+8*4], grid[10+8*4], grid[16+8*4], grid[17+8*4], grid[18+8*4], grid[41]);
   evolve8 e2_10 (grid_evolve[42], grid[1+8*4], grid[2+8*4], grid[3+8*4], grid[9+8*4], grid[11+8*4], grid[17+8*4], grid[18+8*4], grid[19+8*4], grid[42]);
   evolve8 e2_11 (grid_evolve[43], grid[2+8*4], grid[3+8*4], grid[4+8*4], grid[10+8*4], grid[12+8*4], grid[18+8*4], grid[19+8*4], grid[20+8*4], grid[43]);
   evolve8 e2_12 (grid_evolve[44], grid[3+8*4], grid[4+8*4], grid[5+8*4], grid[11+8*4], grid[13+8*4], grid[19+8*4], grid[20+8*4], grid[21+8*4], grid[44]);
   evolve8 e2_13 (grid_evolve[45], grid[4+8*4], grid[5+8*4], grid[6+8*4], grid[12+8*4], grid[14+8*4], grid[20+8*4], grid[21+8*4], grid[22+8*4], grid[45]);
   evolve8 e2_14 (grid_evolve[46], grid[5+8*4], grid[6+8*4], grid[7+8*4], grid[13+8*4], grid[15+8*4], grid[21+8*4], grid[22+8*4], grid[23+8*4], grid[46]);
   evolve5 e2_15 (grid_evolve[47], grid[6+8*4], grid[7+8*4], grid[14+8*4], grid[22+8*4], grid[23+8*4], grid[47]);
    

   evolve5 e6_0 (grid_evolve[48], grid[0+8*5], grid[1+8*5], grid[9+8*5], grid[16+8*5], grid[17+8*5], grid[48]);
   evolve8 e6_1 (grid_evolve[49], grid[0+8*5], grid[1+8*5], grid[2+8*5], grid[8+8*5], grid[10+8*5], grid[16+8*5], grid[17+8*5], grid[18+8*5], grid[49]);
   evolve8 e6_2 (grid_evolve[50], grid[1+8*5], grid[2+8*5], grid[3+8*5], grid[9+8*5], grid[11+8*5], grid[17+8*5], grid[18+8*5], grid[19+8*5], grid[50]);
   evolve8 e6_3 (grid_evolve[51], grid[2+8*5], grid[3+8*5], grid[4+8*5], grid[10+8*5], grid[12+8*5], grid[18+8*5], grid[19+8*5], grid[20+8*5], grid[51]);
   evolve8 e6_4 (grid_evolve[52], grid[3+8*5], grid[4+8*5], grid[5+8*5], grid[11+8*5], grid[13+8*5], grid[19+8*5], grid[20+8*5], grid[21+8*5], grid[52]);
   evolve8 e6_5 (grid_evolve[53], grid[4+8*5], grid[5+8*5], grid[6+8*5], grid[12+8*5], grid[14+8*5], grid[20+8*5], grid[21+8*5], grid[22+8*5], grid[53]);
   evolve8 e6_6 (grid_evolve[54], grid[5+8*5], grid[6+8*5], grid[7+8*5], grid[13+8*5], grid[15+8*5], grid[21+8*5], grid[22+8*5], grid[23+8*5], grid[54]);
   evolve8 e6_7 (grid_evolve[55], grid[6+8*5], grid[7+8*5], grid[48], grid[14+8*5], grid[56], grid[22+8*5], grid[23+8*5], grid[64], grid[47]);
   evolve8 e7_0 (grid_evolve[56], grid[47], grid[0+8*6], grid[1+8*6], grid[55], grid[9+8*6], grid[63], grid[64], grid[65], grid[56]);
   evolve8 e7_1 (grid_evolve[57], grid[0+8*6], grid[1+8*6], grid[2+8*6], grid[8+8*6], grid[10+8*6], grid[64], grid[65], grid[66], grid[57]);
   evolve8 e7_2 (grid_evolve[58], grid[1+8*6], grid[2+8*6], grid[3+8*6], grid[9+8*6], grid[11+8*6], grid[65], grid[66], grid[67], grid[58]);
   evolve8 e7_3 (grid_evolve[59], grid[2+8*6], grid[3+8*6], grid[4+8*6], grid[10+8*6], grid[12+8*6], grid[66], grid[67], grid[68], grid[59]);
   evolve8 e7_4 (grid_evolve[60], grid[3+8*6], grid[4+8*6], grid[5+8*6], grid[11+8*6], grid[13+8*6], grid[67], grid[68], grid[69], grid[60]);
   evolve8 e7_5 (grid_evolve[61], grid[4+8*6], grid[5+8*6], grid[6+8*6], grid[12+8*6], grid[14+8*6], grid[68], grid[69], grid[70], grid[61]);
   evolve8 e7_6 (grid_evolve[62], grid[5+8*6], grid[6+8*6], grid[7+8*6], grid[13+8*6], grid[15+8*6], grid[62]);
   evolve3 e7_7 (grid_evolve[63], grid[6+8*6], grid[7+8*6], grid[14+8*6], grid[63]);
     

   evolve3 e8_0 (grid_evolve[64], grid[0+8*7], grid[1+8*7], grid[9+8*7], grid[0+8*8]);
   evolve5 e8_1 (grid_evolve[65], grid[0+8*7], grid[1+8*7], grid[2+8*7], grid[8+8*7], grid[10+8*7], grid[0+8*8], grid[1+8*8], grid[2+8*8], grid[65]);
   evolve5 e8_2 (grid_evolve[66], grid[1+8*7], grid[2+8*7], grid[3+8*7], grid[9+8*7], grid[11+8*7], grid[1+8*8], grid[2+8*8], grid[3+8*8], grid[66]);
   evolve5 e8_3 (grid_evolve[67], grid[2+8*7], grid[3+8*7], grid[4+8*7], grid[10+8*7], grid[12+8*7], grid[2+8*8], grid[3+8*8], grid[4+8*8], grid[67]);
   evolve5 e8_4 (grid_evolve[68], grid[3+8*7], grid[4+8*7], grid[5+8*7], grid[11+8*7], grid[13+8*7], grid[3+8*8], grid[4+8*8], grid[5+8*8], grid[68]);
   evolve5 e8_5 (grid_evolve[69], grid[4+8*7], grid[5+8*7], grid[6+8*7], grid[12+8*7], grid[14+8*7], grid[4+8*8], grid[5+8*8], grid[6+8*8], grid[69]);
   evolve5 e8_6 (grid_evolve[70], grid[5+8*7], grid[6+8*7], grid[7+8*7], grid[13+8*7], grid[15+8*7], grid[5+8*8], grid[6+8*8], grid[7+8*8], grid[70]);
   evolve3 e8_7 (grid_evolve[71], grid[6+8*7], grid[7+8*7], grid[14+8*7], grid[7+8*8]);

   evolve5 e9_0 (grid_evolve[72], grid[0+8*8], grid[1+8*8], grid[9+8*8], grid[0+8*9], grid[1+8*9], grid[8+8*8], grid[9+8*8], grid[16+8*8], grid[72]);
   evolve8 e9_1 (grid_evolve[73], grid[0+8*8], grid[1+8*8], grid[2+8*8], grid[8+8*8], grid[10+8*8], grid[16+8*8], grid[17+8*8], grid[18+8*8], grid[73]);
   evolve8 e9_2 (grid_evolve[74], grid[1+8*8], grid[2+8*8], grid[3+8*8], grid[9+8*8], grid[11+8*8], grid[17+8*8], grid[18+8*8], grid[19+8*8], grid[74]);
   evolve8 e9_3 (grid_evolve[75], grid[2+8*8], grid[3+8*8], grid[4+8*8], grid[10+8*8], grid[12+8*8], grid[18+8*8], grid[19+8*8], grid[20+8*8], grid[75]);
   evolve8 e9_4 (grid_evolve[76], grid[3+8*8], grid[4+8*8], grid[5+8*8], grid[11+8*8], grid[13+8*8], grid[19+8*8], grid[20+8*8], grid[21+8*8], grid[76]);
   evolve8 e9_5 (grid_evolve[77], grid[4+8*8], grid[5+8*8], grid[6+8*8], grid[12+8*8], grid[14+8*8], grid[20+8*8], grid[21+8*8], grid[22+8*8], grid[77]);
   evolve8 e9_6 (grid_evolve[78], grid[5+8*8], grid[6+8*8], grid[7+8*8], grid[13+8*8], grid[15+8*8], grid[21+8*8], grid[22+8*8], grid[23+8*8], grid[78]);
   evolve5 e9_7 (grid_evolve[79], grid[6+8*8], grid[7+8*8], grid[14+8*8], grid[22+8*8], grid[23+8*8], grid[79]);

   evolve5 e10_0 (grid_evolve[80], grid[0+8*9], grid[1+8*9], grid[9+8*9], grid[0+8*10], grid[1+8*10], grid[8+8*9], grid[9+8*9], grid[16+8*9], grid[80]);
   evolve8 e10_1 (grid_evolve[81], grid[0+8*9], grid[1+8*9], grid[2+8*9], grid[8+8*9], grid[10+8*9], grid[16+8*9], grid[17+8*9], grid[18+8*9], grid[81]);
   evolve8 e10_2 (grid_evolve[82], grid[1+8*9], grid[2+8*9], grid[3+8*9], grid[9+8*9], grid[11+8*9], grid[17+8*9], grid[18+8*9], grid[19+8*9], grid[82]);
   evolve8 e10_3 (grid_evolve[83], grid[2+8*9], grid[3+8*9], grid[4+8*9], grid[10+8*9], grid[12+8*9], grid[18+8*9], grid[19+8*9], grid[20+8*9], grid[83]);
   evolve8 e10_4 (grid_evolve[84], grid[3+8*9], grid[4+8*9], grid[5+8*9], grid[11+8*9], grid[13+8*9], grid[19+8*9], grid[20+8*9], grid[21+8*9], grid[84]);
   evolve8 e10_5 (grid_evolve[85], grid[4+8*9], grid[5+8*9], grid[6+8*9], grid[12+8*9], grid[14+8*9], grid[20+8*9], grid[21+8*9], grid[22+8*9], grid[85]);
   evolve8 e10_6 (grid_evolve[86], grid[5+8*9], grid[6+8*9], grid[7+8*9], grid[13+8*9], grid[15+8*9], grid[21+8*9], grid[22+8*9], grid[23+8*9], grid[86]);
   evolve5 e10_7 (grid_evolve[87], grid[6+8*9], grid[7+8*9], grid[14+8*9], grid[22+8*9], grid[23+8*9], grid[87]);

   evolve5 e11_0 (grid_evolve[88], grid[0+8*10], grid[1+8*10], grid[9+8*10], grid[0+8*11], grid[1+8*11], grid[8+8*10], grid[9+8*10], grid[16+8*10], grid[88]);
   evolve8 e11_1 (grid_evolve[89], grid[0+8*10], grid[1+8*10], grid[2+8*10], grid[8+8*10], grid[10+8*10], grid[16+8*10], grid[17+8*10], grid[18+8*10], grid[89]);
   evolve8 e11_2 (grid_evolve[90], grid[1+8*10], grid[2+8*10], grid[3+8*10], grid[9+8*10], grid[11+8*10], grid[17+8*10], grid[18+8*10], grid[19+8*10], grid[90]);
   evolve8 e11_3 (grid_evolve[91], grid[2+8*10], grid[3+8*10], grid[4+8*10], grid[10+8*10], grid[12+8*10], grid[18+8*10], grid[19+8*10], grid[20+8*10], grid[91]);
   evolve8 e11_4 (grid_evolve[92], grid[3+8*10], grid[4+8*10], grid[5+8*10], grid[11+8*10], grid[13+8*10], grid[19+8*10], grid[20+8*10], grid[21+8*10], grid[92]);
   evolve8 e11_5 (grid_evolve[93], grid[4+8*10], grid[5+8*10], grid[6+8*10], grid[12+8*10], grid[14+8*10], grid[20+8*10], grid[21+8*10], grid[22+8*10], grid[93]);
   evolve8 e11_6 (grid_evolve[94], grid[5+8*10], grid[6+8*10], grid[7+8*10], grid[13+8*10], grid[15+8*10], grid[21+8*10], grid[22+8*10], grid[23+8*10], grid[94]);
   evolve5 e11_7 (grid_evolve[95], grid[6+8*10], grid[7+8*10], grid[14+8*10], grid[22+8*10], grid[23+8*10], grid[95]);

   evolve5 e12_0 (grid_evolve[96], grid[0+8*11], grid[1+8*11], grid[9+8*11], grid[0+8*12], grid[1+8*12], grid[8+8*11], grid[9+8*11], grid[16+8*11], grid[96]);
   evolve8 e12_1 (grid_evolve[97], grid[0+8*11], grid[1+8*11], grid[2+8*11], grid[8+8*11], grid[10+8*11], grid[16+8*11], grid[17+8*11], grid[18+8*11], grid[97]);
   evolve8 e12_2 (grid_evolve[98], grid[1+8*11], grid[2+8*11], grid[3+8*11], grid[9+8*11], grid[11+8*11], grid[17+8*11], grid[18+8*11], grid[19+8*11], grid[98]);
   evolve8 e12_3 (grid_evolve[99], grid[2+8*11], grid[3+8*11], grid[4+8*11], grid[10+8*11], grid[12+8*11], grid[18+8*11], grid[19+8*11], grid[20+8*11], grid[99]);
   evolve8 e12_4 (grid_evolve[100], grid[3+8*11], grid[4+8*11], grid[5+8*11], grid[11+8*11], grid[13+8*11], grid[19+8*11], grid[20+8*11], grid[21+8*11], grid[100]);
   evolve8 e12_5 (grid_evolve[101], grid[4+8*11], grid[5+8*11], grid[6+8*11], grid[12+8*11], grid[14+8*11], grid[20+8*11], grid[21+8*11], grid[22+8*11], grid[101]);
   evolve8 e12_6 (grid_evolve[102], grid[5+8*11], grid[6+8*11], grid[7+8*11], grid[13+8*11], grid[15+8*11], grid[21+8*11], grid[22+8*11], grid[23+8*11]);
   evolve8 e12_7 (grid_evolve[103], grid[6+8*11], grid[7+8*11], grid[14+8*11], grid[22+8*11], grid[23+8*11], grid[103]);

   evolve3 e13_0 (grid_evolve[104], grid[0+8*12], grid[1+8*12], grid[9+8*12], grid[0+8*13]);
   evolve5 e13_1 (grid_evolve[105], grid[0+8*12], grid[1+8*12], grid[2+8*12], grid[8+8*12], grid[10+8*12], grid[9+8*12], grid[16+8*12], grid[17+8*12], grid[105]);
   evolve5 e13_2 (grid_evolve[106], grid[1+8*12], grid[2+8*12], grid[3+8*12], grid[9+8*12], grid[11+8*12], grid[10+8*12], grid[17+8*12], grid[18+8*12], grid[106]);
   evolve5 e13_3 (grid_evolve[107], grid[2+8*12], grid[3+8*12], grid[4+8*12], grid[10+8*12], grid[12+8*12], grid[11+8*12], grid[18+8*12], grid[19+8*12], grid[107]);
   evolve5 e13_4 (grid_evolve[108], grid[3+8*12], grid[4+8*12], grid[5+8*12], grid[11+8*12], grid[13+8*12], grid[12+8*12], grid[19+8*12], grid[20+8*12], grid[108]);
   evolve5 e13_5 (grid_evolve[109], grid[4+8*12], grid[5+8*12], grid[6+8*12], grid[12+8*12], grid[14+8*12], grid[13+8*12], grid[20+8*12], grid[21+8*12], grid[109]);
   evolve5 e13_6 (grid_evolve[110], grid[5+8*12], grid[6+8*12], grid[7+8*12], grid[13+8*12], grid[15+8*12], grid[14+8*12], grid[21+8*12], grid[22+8*12], grid[110]);
   evolve3 e13_7 (grid_evolve[111], grid[6+8*12], grid[7+8*12], grid[14+8*12], grid[111]);

   evolve3 e14_0 (grid_evolve[112], grid[0+8*13], grid[1+8*13], grid[9+8*13], grid[0+8*14]);
   evolve5 e14_1 (grid_evolve[113], grid[0+8*13], grid[1+8*13], grid[2+8*13], grid[8+8*13], grid[10+8*13], grid[9+8*13], grid[16+8*13], grid[17+8*13], grid[113]);
   evolve5 e14_2 (grid_evolve[114], grid[1+8*13], grid[2+8*13], grid[3+8*13], grid[9+8*13], grid[11+8*13], grid[10+8*13], grid[17+8*13], grid[18+8*13], grid[114]);
   evolve5 e14_3 (grid_evolve[115], grid[2+8*13], grid[3+8*13], grid[4+8*13], grid[10+8*13], grid[12+8*13], grid[11+8*13], grid[18+8*13], grid[19+8*13], grid[115]);
   evolve5 e14_4 (grid_evolve[116], grid[3+8*13], grid[4+8*13], grid[5+8*13], grid[11+8*13], grid[13+8*13], grid[12+8*13], grid[19+8*13], grid[20+8*13], grid[116]);
   evolve5 e14_5 (grid_evolve[117], grid[4+8*13], grid[5+8*13], grid[6+8*13], grid[12+8*13], grid[14+8*13], grid[13+8*13], grid[20+8*13], grid[21+8*13], grid[117]);
   evolve5 e14_6 (grid_evolve[118], grid[5+8*13], grid[6+8*13], grid[7+8*13], grid[13+8*13], grid[15+8*13], grid[14+8*13], grid[21+8*13], grid[22+8*13], grid[118]);
   evolve3 e14_7 (grid_evolve[119], grid[6+8*13], grid[7+8*13], grid[14+8*13], grid[119]);

   evolve5 e15_8 (grid_evolve[128], grid[0+8*15], grid[1+8*15], grid[9+8*15], grid[16+8*15], grid[17+8*15], grid[128]);
   evolve8 e15_9 (grid_evolve[129], grid[0+8*15], grid[1+8*15], grid[2+8*15], grid[8+8*15], grid[10+8*15], grid[16+8*15], grid[17+8*15], grid[18+8*15], grid[129]);
   evolve8 e15_10 (grid_evolve[130], grid[1+8*15], grid[2+8*15], grid[3+8*15], grid[9+8*15], grid[11+8*15], grid[17+8*15], grid[18+8*15], grid[19+8*15], grid[130]);
   evolve8 e15_11 (grid_evolve[131], grid[2+8*15], grid[3+8*15], grid[4+8*15], grid[10+8*15], grid[12+8*15], grid[18+8*15], grid[19+8*15], grid[20+8*15], grid[131]);
   evolve8 e15_12 (grid_evolve[132], grid[3+8*15], grid[4+8*15], grid[5+8*15], grid[11+8*15], grid[13+8*15], grid[19+8*15], grid[20+8*15], grid[21+8*15], grid[132]);
   evolve8 e15_13 (grid_evolve[133], grid[4+8*15], grid[5+8*15], grid[6+8*15], grid[12+8*15], grid[14+8*15], grid[20+8*15], grid[21+8*15], grid[22+8*15], grid[133]);
   evolve8 e15_14 (grid_evolve[134], grid[5+8*15], grid[6+8*15], grid[7+8*15], grid[13+8*15], grid[15+8*15], grid[21+8*15], grid[22+8*15], grid[23+8*15], grid[134]);
   evolve5 e15_15 (grid_evolve[135], grid[6+8*15], grid[7+8*15], grid[14+8*15], grid[22+8*15], grid[23+8*15], grid[135]);

   evolve5 e16_0 (grid_evolve[128], grid[0+8*16], grid[1+8*16], grid[9+8*16], grid[16+8*16], grid[17+8*16], grid[128]);
   evolve8 e16_1 (grid_evolve[129], grid[0+8*16], grid[1+8*16], grid[2+8*16], grid[8+8*16], grid[10+8*16], grid[16+8*16], grid[17+8*16], grid[18+8*16], grid[129]);
   evolve8 e16_2 (grid_evolve[130], grid[1+8*16], grid[2+8*16], grid[3+8*16], grid[9+8*16], grid[11+8*16], grid[17+8*16], grid[18+8*16], grid[19+8*16], grid[130]);
   evolve8 e16_3 (grid_evolve[131], grid[2+8*16], grid[3+8*16], grid[4+8*16], grid[10+8*16], grid[12+8*16], grid[18+8*16], grid[19+8*16], grid[20+8*16], grid[131]);
   evolve8 e16_4 (grid_evolve[132], grid[3+8*16], grid[4+8*16], grid[5+8*16], grid[11+8*16], grid[13+8*16], grid[19+8*16], grid[20+8*16], grid[21+8*16], grid[132]);
   evolve8 e16_5 (grid_evolve[133], grid[4+8*16], grid[5+8*16], grid[6+8*16], grid[12+8*16], grid[14+8*16], grid[20+8*16], grid[21+8*16], grid[22+8*16], grid[133]);
   evolve8 e16_6 (grid_evolve[134], grid[5+8*16], grid[6+8*16], grid[7+8*16], grid[13+8*16], grid[15+8*16], grid[21+8*16], grid[22+8*16], grid[23+8*16], grid[134]);
   evolve5 e16_7 (grid_evolve[135], grid[6+8*16], grid[7+8*16], grid[14+8*16], grid[22+8*16], grid[23+8*16], grid[135]);

   evolve5 e17_0 (grid_evolve[136], grid[0+8*17], grid[1+8*17], grid[9+8*17], grid[16+8*17], grid[17+8*17], grid[136]);
   evolve8 e17_1 (grid_evolve[137], grid[0+8*17], grid[1+8*17], grid[2+8*17], grid[8+8*17], grid[10+8*17], grid[16+8*17], grid[17+8*17], grid[18+8*17], grid[137]);
   evolve8 e17_2 (grid_evolve[138], grid[1+8*17], grid[2+8*17], grid[3+8*17], grid[9+8*17], grid[11+8*17], grid[17+8*17], grid[18+8*17], grid[19+8*17], grid[138]);
   evolve8 e17_3 (grid_evolve[139], grid[2+8*17], grid[3+8*17], grid[4+8*17], grid[10+8*17], grid[12+8*17], grid[18+8*17], grid[19+8*17], grid[20+8*17], grid[139]);
   evolve8 e17_4 (grid_evolve[140], grid[3+8*17], grid[4+8*17], grid[5+8*17], grid[11+8*17], grid[13+8*17], grid[19+8*17], grid[20+8*17], grid[21+8*17], grid[140]);
   evolve8 e17_5 (grid_evolve[141], grid[4+8*17], grid[5+8*17], grid[6+8*17], grid[12+8*17], grid[14+8*17], grid[20+8*17], grid[21+8*17], grid[22+8*17], grid[141]);
   evolve8 e17_6 (grid_evolve[142], grid[5+8*17], grid[6+8*17], grid[7+8*17], grid[13+8*17], grid[15+8*17], grid[21+8*17], grid[22+8*17], grid[23+8*17], grid[142]);
   evolve5 e17_7 (grid_evolve[143], grid[6+8*17], grid[7+8*17], grid[14+8*17], grid[22+8*17], grid[23+8*17], grid[143]);

   evolve5 e18_0 (grid_evolve[144], grid[0+8*18], grid[1+8*18], grid[9+8*18], grid[16+8*18], grid[17+8*18], grid[144]);
   evolve8 e18_1 (grid_evolve[145], grid[0+8*18], grid[1+8*18], grid[2+8*18], grid[8+8*18], grid[10+8*18], grid[16+8*18], grid[17+8*18], grid[18+8*18], grid[145]);
   evolve8 e18_2 (grid_evolve[146], grid[1+8*18], grid[2+8*18], grid[3+8*18], grid[9+8*18], grid[11+8*18], grid[17+8*18], grid[18+8*18], grid[19+8*18], grid[146]);
   evolve8 e18_3 (grid_evolve[147], grid[2+8*18], grid[3+8*18], grid[4+8*18], grid[10+8*18], grid[12+8*18], grid[18+8*18], grid[19+8*18], grid[20+8*18], grid[147]);
   evolve8 e18_4 (grid_evolve[148], grid[3+8*18], grid[4+8*18], grid[5+8*18], grid[11+8*18], grid[13+8*18], grid[19+8*18], grid[20+8*18], grid[21+8*18], grid[148]);
   evolve8 e18_5 (grid_evolve[149], grid[4+8*18], grid[5+8*18], grid[6+8*18], grid[12+8*18], grid[14+8*18], grid[20+8*18], grid[21+8*18], grid[22+8*18], grid[149]);
   evolve8 e18_6 (grid_evolve[150], grid[5+8*18], grid[6+8*18], grid[7+8*18], grid[13+8*18], grid[15+8*18], grid[21+8*18], grid[22+8*18], grid[23+8*18], grid[150]);
   evolve5 e18_7 (grid_evolve[151], grid[6+8*18], grid[7+8*18], grid[14+8*18], grid[22+8*18], grid[23+8*18], grid[151]);

   evolve5 e19_0 (grid_evolve[152], grid[0+8*19], grid[1+8*19], grid[9+8*19], grid[16+8*19], grid[17+8*19], grid[152]);
   evolve8 e19_1 (grid_evolve[153], grid[0+8*19], grid[1+8*19], grid[2+8*19], grid[8+8*19], grid[10+8*19], grid[16+8*19], grid[17+8*19], grid[18+8*19], grid[153]);
   evolve8 e19_2 (grid_evolve[154], grid[1+8*19], grid[2+8*19], grid[3+8*19], grid[9+8*19], grid[11+8*19], grid[17+8*19], grid[18+8*19], grid[19+8*19], grid[154]);
   evolve8 e19_3 (grid_evolve[155], grid[2+8*19], grid[3+8*19], grid[4+8*19], grid[10+8*19], grid[12+8*19], grid[18+8*19], grid[19+8*19], grid[20+8*19], grid[155]);
   evolve8 e19_4 (grid_evolve[156], grid[3+8*19], grid[4+8*19], grid[5+8*19], grid[11+8*19], grid[13+8*19], grid[19+8*19], grid[20+8*19], grid[21+8*19], grid[156]);
   evolve8 e19_5 (grid_evolve[157], grid[4+8*19], grid[5+8*19], grid[6+8*19], grid[12+8*19], grid[14+8*19], grid[20+8*19], grid[21+8*19], grid[22+8*19], grid[157]);
   evolve8 e19_6 (grid_evolve[158], grid[5+8*19], grid[6+8*19], grid[7+8*19], grid[13+8*19], grid[15+8*19], grid[21+8*19], grid[22+8*19], grid[23+8*19], grid[158]);
   evolve5 e19_7 (grid_evolve[159], grid[6+8*19], grid[7+8*19], grid[14+8*19], grid[22+8*19], grid[23+8*19], grid[159]);

   evolve3 e20_0 (grid_evolve[160], grid[0+8*20], grid[1+8*20], grid[9+8*20], grid[160]);
   evolve5 e20_1 (grid_evolve[161], grid[0+8*20], grid[1+8*20], grid[2+8*20], grid[8+8*20], grid[10+8*20], grid[161]);
   evolve5 e20_2 (grid_evolve[162], grid[1+8*20], grid[2+8*20], grid[3+8*20], grid[9+8*20], grid[11+8*20], grid[162]);
   evolve5 e20_3 (grid_evolve[163], grid[2+8*20], grid[3+8*20], grid[4+8*20], grid[10+8*20], grid[12+8*20], grid[163]);
   evolve5 e20_4 (grid_evolve[164], grid[3+8*20], grid[4+8*20], grid[5+8*20], grid[11+8*20], grid[13+8*20], grid[164]);
   evolve5 e20_5 (grid_evolve[165], grid[4+8*20], grid[5+8*20], grid[6+8*20], grid[12+8*20], grid[14+8*20], grid[165]);
   evolve5 e20_6 (grid_evolve[166], grid[5+8*20], grid[6+8*20], grid[7+8*20], grid[13+8*20], grid[15+8*20], grid[166]);
   evolve3 e20_7 (grid_evolve[167], grid[6+8*20], grid[7+8*20], grid[14+8*20], grid[167]);

   evolve5 e21_0 (grid_evolve[168], grid[0+8*21], grid[1+8*21], grid[9+8*21], grid[160+8*1], grid[161+8*1], grid[168]);
   evolve8 e21_1 (grid_evolve[169], grid[0+8*21], grid[1+8*21], grid[2+8*21], grid[8+8*21], grid[10+8*21], grid[160+8*1], grid[161+8*1], grid[162+8*1], grid[169]);
   evolve8 e21_2 (grid_evolve[170], grid[1+8*21], grid[2+8*21], grid[3+8*21], grid[9+8*21], grid[11+8*21], grid[161+8*1], grid[162+8*1], grid[163+8*1], grid[170]);
   evolve8 e21_3 (grid_evolve[171], grid[2+8*21], grid[3+8*21], grid[4+8*21], grid[10+8*21], grid[12+8*21], grid[162+8*1], grid[163+8*1], grid[164+8*1], grid[171]);
   evolve8 e21_4 (grid_evolve[172], grid[3+8*21], grid[4+8*21], grid[5+8*21], grid[11+8*21], grid[13+8*21], grid[163+8*1], grid[164+8*1], grid[165+8*1], grid[172]);
   evolve8 e21_5 (grid_evolve[173], grid[4+8*21], grid[5+8*21], grid[6+8*21], grid[12+8*21], grid[14+8*21], grid[164+8*1], grid[165+8*1], grid[166+8*1], grid[173]);
   evolve8 e21_6 (grid_evolve[174], grid[5+8*21], grid[6+8*21], grid[7+8*21], grid[13+8*21], grid[15+8*21], grid[165+8*1], grid[166+8*1], grid[167+8*1], grid[174]);
   evolve5 e21_7 (grid_evolve[175], grid[6+8*21], grid[7+8*21], grid[14+8*21], grid[166+8*1], grid[167+8*1], grid[175]);

   evolve3 e22_0 (grid_evolve[176], grid[0+8*22], grid[1+8*22], grid[9+8*22], grid[176]);
   evolve5 e22_1 (grid_evolve[177], grid[0+8*22], grid[1+8*22], grid[2+8*22], grid[8+8*22], grid[10+8*22], grid[177]);
   evolve5 e22_2 (grid_evolve[178], grid[1+8*22], grid[2+8*22], grid[3+8*22], grid[9+8*22], grid[11+8*22], grid[178]);
   evolve5 e22_3 (grid_evolve[179], grid[2+8*22], grid[3+8*22], grid[4+8*22], grid[10+8*22], grid[12+8*22], grid[179]);
   evolve5 e22_4 (grid_evolve[180], grid[3+8*22], grid[4+8*22], grid[5+8*22], grid[11+8*22], grid[13+8*22], grid[180]);
   evolve5 e22_5 (grid_evolve[181], grid[4+8*22], grid[5+8*22], grid[6+8*22], grid[12+8*22], grid[14+8*22], grid[181]);
   evolve5 e22_6 (grid_evolve[182], grid[5+8*22], grid[6+8*22], grid[7+8*22], grid[13+8*22], grid[15+8*22], grid[182]);
   evolve3 e22_7 (grid_evolve[183], grid[6+8*22], grid[7+8*22], grid[14+8*22], grid[183]);

   evolve5 e23_0 (grid_evolve[184], grid[0+8*23], grid[1+8*23], grid[9+8*23], grid[176+8*1], grid[177+8*1], grid[184]);
   evolve8 e23_1 (grid_evolve[185], grid[0+8*23], grid[1+8*23], grid[2+8*23], grid[8+8*23], grid[10+8*23], grid[176+8*1], grid[177+8*1], grid[178+8*1], grid[185]);
   evolve8 e23_2 (grid_evolve[186], grid[1+8*23], grid[2+8*23], grid[3+8*23], grid[9+8*23], grid[11+8*23], grid[177+8*1], grid[178+8*1], grid[179+8*1], grid[186]);
   evolve8 e23_3 (grid_evolve[187], grid[2+8*23], grid[3+8*23], grid[4+8*23], grid[10+8*23], grid[12+8*23], grid[178+8*1], grid[179+8*1], grid[180+8*1], grid[187]);
   evolve8 e23_4 (grid_evolve[188], grid[3+8*23], grid[4+8*23], grid[5+8*23], grid[11+8*23], grid[13+8*23], grid[179+8*1], grid[180+8*1], grid[181+8*1], grid[188]);
   evolve8 e23_5 (grid_evolve[189], grid[4+8*23], grid[5+8*23], grid[6+8*23], grid[12+8*23], grid[14+8*23], grid[180+8*1], grid[181+8*1], grid[182+8*1], grid[189]);
   evolve8 e23_6 (grid_evolve[190], grid[5+8*23], grid[6+8*23], grid[7+8*23], grid[13+8*23], grid[15+8*23], grid[181+8*1], grid[182+8*1], grid[183+8*1], grid[190]);
   evolve5 e23_7 (grid_evolve[191], grid[6+8*23], grid[7+8*23], grid[14+8*23], grid[182+8*1], grid[183+8*1], grid[191]);

   evolve3 e24_0 (grid_evolve[192], grid[0+8*24], grid[1+8*24], grid[9+8*24], grid[192]);
   evolve5 e24_1 (grid_evolve[193], grid[0+8*24], grid[1+8*24], grid[2+8*24], grid[8+8*24], grid[10+8*24], grid[193]);
   evolve5 e24_2 (grid_evolve[194], grid[1+8*24], grid[2+8*24], grid[3+8*24], grid[9+8*24], grid[11+8*24], grid[194]);
   evolve5 e24_3 (grid_evolve[195], grid[2+8*24], grid[3+8*24], grid[4+8*24], grid[10+8*24], grid[12+8*24], grid[195]);
   evolve5 e24_4 (grid_evolve[196], grid[3+8*24], grid[4+8*24], grid[5+8*24], grid[11+8*24], grid[13+8*24], grid[196]);
   evolve5 e24_5 (grid_evolve[197], grid[4+8*24], grid[5+8*24], grid[6+8*24], grid[12+8*24], grid[14+8*24], grid[197]);
   evolve5 e24_6 (grid_evolve[198], grid[5+8*24], grid[6+8*24], grid[7+8*24], grid[13+8*24], grid[15+8*24], grid[198]);
   evolve3 e24_7 (grid_evolve[199], grid[6+8*24], grid[7+8*24], grid[14+8*24], grid[199]);

   evolve5 e25_0 (grid_evolve[200], grid[0+8*25], grid[1+8*25], grid[9+8*25], grid[16+8*25], grid[17+8*25], grid[200]);
   evolve8 e25_1 (grid_evolve[201], grid[0+8*25], grid[1+8*25], grid[2+8*25], grid[8+8*25], grid[10+8*25], grid[16+8*25], grid[17+8*25], grid[18+8*25], grid[201]);
   evolve8 e25_2 (grid_evolve[202], grid[1+8*25], grid[2+8*25], grid[3+8*25], grid[9+8*25], grid[11+8*25], grid[17+8*25], grid[18+8*25], grid[19+8*25], grid[202]);
   evolve8 e25_3 (grid_evolve[203], grid[2+8*25], grid[3+8*25], grid[4+8*25], grid[10+8*25], grid[12+8*25], grid[18+8*25], grid[19+8*25], grid[20+8*25], grid[203]);
   evolve8 e25_4 (grid_evolve[204], grid[3+8*25], grid[4+8*25], grid[5+8*25], grid[11+8*25], grid[13+8*25], grid[19+8*25], grid[20+8*25], grid[21+8*25], grid[204]);
   evolve8 e25_5 (grid_evolve[205], grid[4+8*25], grid[5+8*25], grid[6+8*25], grid[12+8*25], grid[14+8*25], grid[20+8*25], grid[21+8*25], grid[22+8*25], grid[205]);
   evolve8 e25_6 (grid_evolve[206], grid[5+8*25], grid[6+8*25], grid[7+8*25], grid[13+8*25], grid[15+8*25], grid[21+8*25], grid[22+8*25], grid[23+8*25], grid[206]);
   evolve5 e25_7 (grid_evolve[207], grid[6+8*25], grid[7+8*25], grid[14+8*25], grid[22+8*25], grid[23+8*25], grid[207]);

   evolve3 e26_0 (grid_evolve[208], grid[0+8*26], grid[1+8*26], grid[9+8*26], grid[208]);
   evolve5 e26_1 (grid_evolve[209], grid[0+8*26], grid[1+8*26], grid[2+8*26], grid[8+8*26], grid[10+8*26], grid[209]);
   evolve5 e26_2 (grid_evolve[210], grid[1+8*26], grid[2+8*26], grid[3+8*26], grid[9+8*26], grid[11+8*26], grid[210]);
   evolve5 e26_3 (grid_evolve[211], grid[2+8*26], grid[3+8*26], grid[4+8*26], grid[10+8*26], grid[12+8*26], grid[211]);
   evolve5 e26_4 (grid_evolve[212], grid[3+8*26], grid[4+8*26], grid[5+8*26], grid[11+8*26], grid[13+8*26], grid[212]);
   evolve5 e26_5 (grid_evolve[213], grid[4+8*26], grid[5+8*26], grid[6+8*26], grid[12+8*26], grid[14+8*26], grid[213]);
   evolve5 e26_6 (grid_evolve[214], grid[5+8*26], grid[6+8*26], grid[7+8*26], grid[13+8*26], grid[15+8*26], grid[214]);
   evolve3 e26_7 (grid_evolve[215], grid[6+8*26], grid[7+8*26], grid[14+8*26], grid[215]);

   evolve5 e27_0 (grid_evolve[216], grid[0+8*27], grid[1+8*27], grid[9+8*27], grid[16+8*27], grid[17+8*27], grid[216]);
   evolve8 e27_1 (grid_evolve[217], grid[0+8*27], grid[1+8*27], grid[2+8*27], grid[8+8*27], grid[10+8*27], grid[16+8*27], grid[17+8*27], grid[18+8*27], grid[217]);
   evolve8 e27_2 (grid_evolve[218], grid[1+8*27], grid[2+8*27], grid[3+8*27], grid[9+8*27], grid[11+8*27], grid[17+8*27], grid[18+8*27], grid[19+8*27], grid[218]);
   evolve8 e27_3 (grid_evolve[219], grid[2+8*27], grid[3+8*27], grid[4+8*27], grid[10+8*27], grid[12+8*27], grid[18+8*27], grid[19+8*27], grid[20+8*27], grid[219]);
   evolve8 e27_4 (grid_evolve[220], grid[3+8*27], grid[4+8*27], grid[5+8*27], grid[11+8*27], grid[13+8*27], grid[19+8*27], grid[20+8*27], grid[21+8*27], grid[220]);
   evolve8 e27_5 (grid_evolve[221], grid[4+8*27], grid[5+8*27], grid[6+8*27], grid[12+8*27], grid[14+8*27], grid[20+8*27], grid[21+8*27], grid[22+8*27], grid[221]);
   evolve8 e27_6 (grid_evolve[222], grid[5+8*27], grid[6+8*27], grid[7+8*27], grid[13+8*27], grid[15+8*27], grid[21+8*27], grid[22+8*27], grid[23+8*27], grid[222]);
   evolve5 e27_7 (grid_evolve[223], grid[6+8*27], grid[7+8*27], grid[14+8*27], grid[22+8*27], grid[23+8*27], grid[223]);

   evolve3 e28_0 (grid_evolve[224], grid[0+8*28], grid[1+8*28], grid[9+8*28], grid[224]);
   evolve5 e28_1 (grid_evolve[225], grid[0+8*28], grid[1+8*28], grid[2+8*28], grid[8+8*28], grid[10+8*28], grid[225]);
   evolve5 e28_2 (grid_evolve[226], grid[1+8*28], grid[2+8*28], grid[3+8*28], grid[9+8*28], grid[11+8*28], grid[226]);
   evolve5 e28_3 (grid_evolve[227], grid[2+8*28], grid[3+8*28], grid[4+8*28], grid[10+8*28], grid[12+8*28], grid[227]);
   evolve5 e28_4 (grid_evolve[228], grid[3+8*28], grid[4+8*28], grid[5+8*28], grid[11+8*28], grid[13+8*28], grid[228]);
   evolve5 e28_5 (grid_evolve[229], grid[4+8*28], grid[5+8*28], grid[6+8*28], grid[12+8*28], grid[14+8*28], grid[229]);
   evolve5 e28_6 (grid_evolve[230], grid[5+8*28], grid[6+8*28], grid[7+8*28], grid[13+8*28], grid[15+8*28], grid[230]);
   evolve3 e28_7 (grid_evolve[231], grid[6+8*28], grid[7+8*28], grid[14+8*28], grid[231]);

   evolve5 e29_0 (grid_evolve[232], grid[0+8*29], grid[1+8*29], grid[9+8*29], grid[16+8*29], grid[17+8*29], grid[232]);
   evolve8 e29_1 (grid_evolve[233], grid[0+8*29], grid[1+8*29], grid[2+8*29], grid[8+8*29], grid[10+8*29], grid[16+8*29], grid[17+8*29], grid[18+8*29], grid[233]);
   evolve8 e29_2 (grid_evolve[234], grid[1+8*29], grid[2+8*29], grid[3+8*29], grid[9+8*29], grid[11+8*29], grid[17+8*29], grid[18+8*29], grid[19+8*29], grid[234]);
   evolve8 e29_3 (grid_evolve[235], grid[2+8*29], grid[3+8*29], grid[4+8*29], grid[10+8*29], grid[12+8*29], grid[18+8*29], grid[19+8*29], grid[20+8*29], grid[235]);
   evolve8 e29_4 (grid_evolve[236], grid[3+8*29], grid[4+8*29], grid[5+8*29], grid[11+8*29], grid[13+8*29], grid[19+8*29], grid[20+8*29], grid[21+8*29], grid[236]);
   evolve8 e29_5 (grid_evolve[237], grid[4+8*29], grid[5+8*29], grid[6+8*29], grid[12+8*29], grid[14+8*29], grid[20+8*29], grid[21+8*29], grid[22+8*29], grid[237]);
   evolve8 e29_6 (grid_evolve[238], grid[5+8*29], grid[6+8*29], grid[7+8*29], grid[13+8*29], grid[15+8*29], grid[21+8*29], grid[22+8*29], grid[23+8*29], grid[238]);
   evolve5 e29_7 (grid_evolve[239], grid[6+8*29], grid[7+8*29], grid[14+8*29], grid[22+8*29], grid[23+8*29], grid[239]);

   evolve5 e30_0 (grid_evolve[240], grid[0+8*30], grid[1+8*30], grid[9+8*30], grid[16+8*30], grid[17+8*30], grid[240]);
   evolve8 e30_1 (grid_evolve[241], grid[0+8*30], grid[1+8*30], grid[2+8*30], grid[8+8*30], grid[10+8*30], grid[16+8*30], grid[17+8*30], grid[18+8*30], grid[241]);
   evolve8 e30_2 (grid_evolve[242], grid[1+8*30], grid[2+8*30], grid[3+8*30], grid[9+8*30], grid[11+8*30], grid[17+8*30], grid[18+8*30], grid[19+8*30], grid[242]);
   evolve8 e30_3 (grid_evolve[243], grid[2+8*30], grid[3+8*30], grid[4+8*30], grid[10+8*30], grid[12+8*30], grid[18+8*30], grid[19+8*30], grid[20+8*30], grid[243]);
   evolve8 e30_4 (grid_evolve[244], grid[3+8*30], grid[4+8*30], grid[5+8*30], grid[11+8*30], grid[13+8*30], grid[19+8*30], grid[20+8*30], grid[21+8*30], grid[244]);
   evolve8 e30_5 (grid_evolve[245], grid[4+8*30], grid[5+8*30], grid[6+8*30], grid[12+8*30], grid[14+8*30], grid[20+8*30], grid[21+8*30], grid[22+8*30], grid[245]);
   evolve8 e30_6 (grid_evolve[246], grid[5+8*30], grid[6+8*30], grid[7+8*30], grid[13+8*30], grid[15+8*30], grid[21+8*30], grid[22+8*30], grid[23+8*30], grid[246]);
   evolve5 e30_7 (grid_evolve[247], grid[6+8*30], grid[7+8*30], grid[14+8*30], grid[22+8*30], grid[23+8*30], grid[247]);

   evolve3 e31_0 (grid_evolve[248], grid[0+8*31], grid[1+8*31], grid[9+8*31], grid[248]);
   evolve5 e31_1 (grid_evolve[249], grid[0+8*31], grid[1+8*31], grid[2+8*31], grid[8+8*31], grid[10+8*31], grid[249]);
   evolve5 e31_2 (grid_evolve[250], grid[1+8*31], grid[2+8*31], grid[3+8*31], grid[9+8*31], grid[11+8*31], grid[250]);
   evolve5 e31_3 (grid_evolve[251], grid[2+8*31], grid[3+8*31], grid[4+8*31], grid[10+8*31], grid[12+8*31], grid[251]);
   evolve5 e31_4 (grid_evolve[252], grid[3+8*31], grid[4+8*31], grid[5+8*31], grid[11+8*31], grid[13+8*31], grid[252]);
   evolve5 e31_5 (grid_evolve[253], grid[4+8*31], grid[5+8*31], grid[6+8*31], grid[12+8*31], grid[14+8*31], grid[253]);
   evolve5 e31_6 (grid_evolve[254], grid[5+8*31], grid[6+8*31], grid[7+8*31], grid[13+8*31], grid[15+8*31], grid[254]);
   evolve3 e31_7 (grid_evolve[255], grid[6+8*31], grid[7+8*31], grid[14+8*31], grid[255]);




 
endmodule // top


module evolve3 (next_state, vector1, vector2, vector3, current_state);
	
   input logic  vector1;
   input logic  vector2;
   input logic  vector3;
   input logic  current_state;
   output logic next_state;
   
   logic [3:0] 	sum;
   
   assign sum = vector1 + vector2 + vector3;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve3

module evolve5 (next_state, vector1, vector2, vector3, 
		vector4, vector5, current_state);
   
   input logic   vector1;
   input logic 	 vector2;
   input logic 	 vector3;
   input logic 	 vector4;
   input logic 	 vector5;
   input logic 	 current_state;
   output logic  next_state;
   
   logic [3:0] 	 sum;
   
   assign sum = vector1 + vector2 + vector3 + vector4 + vector5;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve5


module evolve8 (next_state, vector1, vector2, vector3, 
		vector4, vector5, vector6, 
		vector7, vector8, current_state);
   
   input logic 	vector1;
   input logic 	vector2;
   input logic 	vector3;
   input logic 	vector4;
   input logic 	vector5;
	
   input logic 	vector6;
   input logic 	vector7;
   input logic 	vector8;
   input logic 	current_state;
   output logic next_state;
   
   logic [3:0] 	sum;
   
   assign sum = vector1 + vector2 + vector3 + vector4 + 
		vector5 + vector6 + vector7 + vector8;
   rules r1 (sum, current_state, next_state);
   
endmodule // evolve8


module rules (pop_count, current_state, next_state);
   
   input logic [3:0] pop_count;
   input logic 	     current_state;
   output logic      next_state;
   
   assign next_state = (pop_count == 2 & current_state) | pop_count == 3;
   
endmodule // rules

module New_Datapath (grid, reset, clk, q);
input logic [255:0] grid;
input logic reset;
input logic clk;
output logic [255:0] q;
logic [255:0] grid_evolve;

FSM sw(clk, reset, en, rst);
mux2 #(256) m1(.d1(grid), .d0(q), .s(rst), .y(outputY));
datapath dp(.grid(outputY), .grid_evolve(grid_evolve));
flopenr #(256)f1 (.clk(clk), .reset(rst), .en(en), .d(grid_evolve), .q(q));



endmodule


